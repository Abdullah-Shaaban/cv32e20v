module xif_sva (
    input  logic clk_i,
    input  logic rst_ni
);


endmodule : xif_sva